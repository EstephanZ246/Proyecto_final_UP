module instancias(/*program_counter*/
                  clk,/*reloj general*/
                  reset_program_counter,/*reset de program_counter*/
                  enable_program__counter,/*enable de program_counter*/
                  load_program_counter,/*entrada para cargar el address_RAM */
                  address_RAM,/*program_counter*/
                  PC,/*program_counter*/


                            );
